----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:27:35 10/09/2017 
-- Design Name: 
-- Module Name:    Mux - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Mux is
    Port ( i : in  STD_LOGIC;
           Crs2 : in  STD_LOGIC_VECTOR (31 downto 0);
           E_seu : in  STD_LOGIC_VECTOR (31 downto 0);
           S_mux : out  STD_LOGIC_VECTOR (31 downto 0));
end Mux;

architecture Behavioral of Mux is

begin

process(i,E_seu,Crs2)
begin
	if(i='1')then
	   S_mux<= E_seu;
	else 
		if(i='0')then
			S_mux <= Crs2;
		end if ; 
end if;

end process;
end Behavioral;

